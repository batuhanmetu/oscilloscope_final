module static2
	(
		input wire clk, 
		output wire [2:0] red,
		output wire [2:0] green,
		output wire [2:0] blue,
		input wire [9:0] x,
		input wire [9:0] y,
		input wire video_on
	);
	
	reg [2:0] rgb_red;
	reg [2:0] rgb_green;
	reg [2:0] rgb_blue;
	

        always @(posedge clk)
		  begin
		  if( x >= 160  )
		  begin
        if( ((x%40==0 && y%2==0) || (x%2==0 && y%40==0)) && y != 240 && x != 160 )
			  begin
				rgb_red <= 3'b111;
				rgb_blue <= 3'b111;
				rgb_green <= 3'b111;
			  end
		  else if ( y==240 || x==160 )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
			else
				begin
				rgb_red <= 3'b000;
				rgb_blue <= 3'b000;
				rgb_green <= 3'b000;
				end			
		 end
		 else if ((y==100 && (x== 10 || x== 11 ||  x== 12)) ||   // V
					 (y==101 && (x== 11 || x== 12 ||  x== 13)) ||   
					 (y==102 && (x== 12 || x== 13 ||  x== 14)) ||
					 (y==103 && (x== 13 || x== 14 ||  x== 15)) ||
					 (y==104 && (x== 14 || x== 15 ||  x== 16)) ||
					 (y==105 && (x== 15 || x== 16 ||  x== 17)) ||
					 (y==106 && (x== 16 || x== 17 ||  x== 18)) ||
					 (y==107 && (x== 17 || x== 18 ||  x== 19)) ||
					 (y==108 && (x== 18 || x== 19 ||  x== 20)) ||
					 (y==109 && (x== 19 || x== 20 ||  x== 21)) ||
					 (y==110 && (x== 20 || x== 21 ||  x== 22)) ||
					 (y==111 && (x== 21 || x== 22 ||  x== 23)) ||
					 (y==110 && (x== 22 || x== 23 ||  x== 24)) ||
					 (y==109 && (x== 23 || x== 24 ||  x== 25)) ||
					 (y==108 && (x== 24 || x== 25 ||  x== 26)) ||
					 (y==107 && (x== 25 || x== 26 ||  x== 27)) ||
					 (y==106 && (x== 26 || x== 27 ||  x== 28)) ||
					 (y==105 && (x== 27 || x== 28 ||  x== 29)) ||
					 (y==104 && (x== 28 || x== 29 ||  x== 30)) ||
					 (y==103 && (x== 29 || x== 30 ||  x== 31)) ||
					 (y==102 && (x== 30 || x== 31 ||  x== 32)) ||
					 (y==101 && (x== 31 || x== 32 ||  x== 33)) ||
					 (y==100 && (x== 32 || x== 33 ||  x== 34)) )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
			else if ( (y > 104 && y < 120) && ( x== 34 || x== 35 ) || // p
					(y==106 && (x== 36 || x== 37 )) ||
					(y==107 && (x== 37 || x== 38 )) ||
					(y==108 && (x== 38 || x== 39 )) ||
					(y==109 && (x== 39 || x== 40 )) ||
					(y==110 && (x== 39 || x== 40 )) ||
					(y==111 && (x== 38 || x== 39 )) ||
					(y==112 && (x== 37 || x== 38 )) ||
					(y==113 && (x== 36 || x== 37 )) )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				else if ( (y > 104 && y < 120) && ( x== 44 || x== 45 ) || // p
					(y==106 && (x== 46 || x== 47 )) ||
					(y==107 && (x== 47 || x== 48 )) ||
					(y==108 && (x== 48 || x== 49 )) ||
					(y==109 && (x== 49 || x== 50 )) ||
					(y==110 && (x== 49 || x== 50 )) ||
					(y==111 && (x== 48 || x== 49 )) ||
					(y==112 && (x== 47 || x== 48 )) ||
					(y==113 && (x== 46 || x== 47 )) )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				else if ( ((y == 104 ) && ( x > 55 && x < 66 ))  ||  			 //=
							 ((y == 108 ) && ( x > 55 && x < 66))   ||
							 ((y == 184 ) && ( x > 55 && x < 66 ))  ||  		
							 ((y == 188 ) && ( x > 55 && x < 66))   ||	
							 ((y == 264 ) && ( x > 55 && x < 66 ))  ||  		
							 ((y == 268 ) && ( x > 55 && x < 66))   ||
							 ((y == 344 ) && ( x > 55 && x < 66 ))  ||  		
							 ((y == 348 ) && ( x > 55 && x < 66))	 )	
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				
				else if ((y==180 && (x== 10 || x== 11 ||  x== 12)) ||   // V
							 (y==181 && (x== 11 || x== 12 ||  x== 13)) ||   
							 (y==182 && (x== 12 || x== 13 ||  x== 14)) ||
							 (y==183 && (x== 13 || x== 14 ||  x== 15)) ||
							 (y==184 && (x== 14 || x== 15 ||  x== 16)) ||
							 (y==185 && (x== 15 || x== 16 ||  x== 17)) ||
							 (y==186 && (x== 16 || x== 17 ||  x== 18)) ||
							 (y==187 && (x== 17 || x== 18 ||  x== 19)) ||
							 (y==188 && (x== 18 || x== 19 ||  x== 20)) ||
							 (y==189 && (x== 19 || x== 20 ||  x== 21)) ||
							 (y==190 && (x== 20 || x== 21 ||  x== 22)) ||
							 (y==191 && (x== 21 || x== 22 ||  x== 23)) ||
							 (y==190 && (x== 22 || x== 23 ||  x== 24)) ||
							 (y==189 && (x== 23 || x== 24 ||  x== 25)) ||
							 (y==188 && (x== 24 || x== 25 ||  x== 26)) ||
							 (y==187 && (x== 25 || x== 26 ||  x== 27)) ||
							 (y==186 && (x== 26 || x== 27 ||  x== 28)) ||
							 (y==185 && (x== 27 || x== 28 ||  x== 29)) ||
							 (y==184 && (x== 28 || x== 29 ||  x== 30)) ||
							 (y==183 && (x== 29 || x== 30 ||  x== 31)) ||
							 (y==182 && (x== 30 || x== 31 ||  x== 32)) ||
							 (y==181 && (x== 31 || x== 32 ||  x== 33)) ||
							 (y==180 && (x== 32 || x== 33 ||  x== 34)) )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				
				else if (                                          //m
							(y==193 && (x== 33 || x== 34 )) ||
							(y==192 && (x== 33 || x== 34 )) ||
							(y==191 && (x== 33 || x== 34 )) ||
							(y==190 && (x== 33 || x== 34 )) ||
							(y==189 && (x== 33 || x== 34 )) ||
							(y==188 && (x== 33 || x== 34 )) ||
							(y==187 && (x== 34 || x== 35 )) ||
							(y==186 && (x== 35 || x== 36 )) ||
							(y==186 && (x== 36 || x== 37 )) ||
							(y==187 && (x== 37 || x== 38 )) ||
							
					
							(y==193 && (x== 38 || x== 39 )) ||
							(y==192 && (x== 38 || x== 39 )) ||
							(y==191 && (x== 38 || x== 39 )) ||
							(y==190 && (x== 38 || x== 39 )) ||
							(y==189 && (x== 38 || x== 39 )) ||
							(y==188 && (x== 38 || x== 39 )) ||
							(y==187 && (x== 39 || x== 40 )) ||
							(y==186 && (x== 40 || x== 41 )) ||
							(y==186 && (x== 41 || x== 42 )) ||
							(y==187 && (x== 42 || x== 43 )) ||
							(y==188 && (x== 43 || x== 44 )) ||
							(y==189 && (x== 43 || x== 44 )) ||
							(y==190 && (x== 43 || x== 44 )) ||
							(y==191 && (x== 43 || x== 44 )) ||
							(y==192 && (x== 43 || x== 44 )) ||
							(y==193 && (x== 43 || x== 44 ))   )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				
				else if  ((y==260 && (x== 0 || x== 1 ||  x== 2)) ||   // V
							 (y==261 && (x== 1 || x== 2 ||  x== 3)) ||   
							 (y==262 && (x== 2 || x== 3 ||  x== 4)) ||
							 (y==263 && (x== 3 || x== 4 ||  x== 5)) ||
							 (y==264 && (x== 4 || x== 5 ||  x== 6)) ||
							 (y==265 && (x== 5 || x== 6 ||  x== 7)) ||
							 (y==266 && (x== 6 || x== 7 ||  x== 8)) ||
							 (y==267 && (x== 7 || x== 8 ||  x== 9)) ||
							 (y==268 && (x== 8 || x== 9 ||  x== 10)) ||
							 (y==269 && (x== 9 || x== 10 ||  x== 11)) ||
							 (y==270 && (x== 10 || x== 11 ||  x== 12)) ||
							 (y==271 && (x== 11 || x== 12 ||  x== 13)) ||
							 (y==270 && (x== 12 || x== 13 ||  x== 14)) ||
							 (y==269 && (x== 13 || x== 14 ||  x== 15)) ||
							 (y==268 && (x== 14 || x== 15 ||  x== 16)) ||
							 (y==267 && (x== 15 || x== 16 ||  x== 17)) ||
							 (y==266 && (x== 16 || x== 17 ||  x== 18)) ||
							 (y==265 && (x== 17 || x== 18 ||  x== 19)) ||
							 (y==264 && (x== 18 || x== 19 ||  x== 20)) ||
							 (y==263 && (x== 19 || x== 20 ||  x== 21)) ||
							 (y==262 && (x== 20 || x== 21 ||  x== 22)) ||
							 (y==261 && (x== 21 || x== 22 ||  x== 23)) ||
							 (y==260 && (x== 22 || x== 23 ||  x== 24)) )
						begin
							rgb_red <= 3'b111;
							rgb_blue <= 3'b111;
							rgb_green <= 3'b111;
						end
					 else if((y==273 && (x== 23 || x== 24 )) ||   		 //r
								(y==272 && (x== 23 || x== 24 )) ||
								(y==271 && (x== 23 || x== 24 )) ||
								(y==270 && (x== 23 || x== 24 )) ||
								(y==269 && (x== 23 || x== 24 )) ||
								(y==268 && (x== 23 || x== 24 )) ||
								(y==267 && (x== 24 || x== 25 )) ||
								(y==266 && (x== 25 || x== 26 )) ||
								(y==266 && (x== 26 || x== 27 )) ||
								(y==267 && (x== 27 || x== 28 )) ||
								(y==267 && (x== 28 || x== 29 )) ||	
								(y==267 && (x== 29 || x== 30 ))	)
					 begin
							rgb_red <= 3'b111;
							rgb_blue <= 3'b111;
							rgb_green <= 3'b111;
					 end
					
					else if (                                          //m
							(y==273 && (x== 33 || x== 34 )) ||
							(y==272 && (x== 33 || x== 34 )) ||
							(y==271 && (x== 33 || x== 34 )) ||
							(y==270 && (x== 33 || x== 34 )) ||
							(y==269 && (x== 33 || x== 34 )) ||
							(y==268 && (x== 33 || x== 34 )) ||
							(y==267 && (x== 34 || x== 35 )) ||
							(y==266 && (x== 35 || x== 36 )) ||
							(y==266 && (x== 36 || x== 37 )) ||
							(y==267 && (x== 37 || x== 38 )) ||
							
					
							(y==273 && (x== 38 || x== 39 )) ||
							(y==272 && (x== 38 || x== 39 )) ||
							(y==271 && (x== 38 || x== 39 )) ||
							(y==270 && (x== 38 || x== 39 )) ||
							(y==269 && (x== 38 || x== 39 )) ||
							(y==268 && (x== 38 || x== 39 )) ||
							(y==267 && (x== 39 || x== 40 )) ||
							(y==266 && (x== 40 || x== 41 )) ||
							(y==266 && (x== 41 || x== 42 )) ||
							(y==267 && (x== 42 || x== 43 )) ||
							(y==268 && (x== 43 || x== 44 )) ||
							(y==269 && (x== 43 || x== 44 )) ||
							(y==270 && (x== 43 || x== 44 )) ||
							(y==271 && (x== 43 || x== 44 )) ||
							(y==272 && (x== 43 || x== 44 )) ||
							(y==273 && (x== 43 || x== 44 ))   )
				begin
					rgb_red <= 3'b111;
					rgb_blue <= 3'b111;
					rgb_green <= 3'b111;
				end
				else if ((y==266 && (x== 49 || x== 50 )) ||      //s
							(y==267 && (x== 48 || x== 51 )) ||
							(y==268 && (x== 48 )) ||
							(y==269 && (x== 49 || x== 50 )) ||
							(y==270 && (x== 51 )) ||
							(y==271 && (x== 48 || x== 51 )) ||
							(y==272 && (x== 49 || x== 50 ))     )	
				begin
						rgb_red <= 3'b111;
						rgb_blue <= 3'b111;
						rgb_green <= 3'b111;
				end	
				
				else if ( ((y==335) && (x==35 || x==36)) ||      //f
							 ((y==336) && (x==34 || x==35 || x==37 || x==38)) ||
							 ((y==337) && (x==33 || x==34 || x==38 || x==39)) ||
							 ((y==338) && (x==32 || x==33 || x==39 || x==40)) ||
							 ((y==339) && (x==31 || x==32 || x==40 || x==41)) ||
							 ((y==340) && (x==30 || x==31 || x==41 || x==42)) ||
							 ((y>=341  && y<= 360) && (x==30 || x==31)) ||
							 ((y==348 || y==349 ) && (x==27||x==28||x==29 || x==30 ||x==31 || x==32 || x==33 || x==34))
							 )
				begin
						rgb_red <= 3'b111;
						rgb_blue <= 3'b111;
						rgb_green <= 3'b111;
				end	

		
        	else 
				begin
				rgb_red <= 3'b000;
				rgb_blue <= 3'b000;
				rgb_green <= 3'b000;
				end
		  
		end
        // output
        assign red = (video_on) ? rgb_red : 3'b0;
		  assign green = (video_on) ? rgb_green : 3'b0;
		  assign blue = (video_on) ? rgb_blue : 3'b0;

endmodule